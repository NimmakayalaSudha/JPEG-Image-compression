`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/20/2021 10:23:56 AM
// Design Name: 
// Module Name: obc_new
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module obc_new(x1,x2,x3,x4,x5,x6,x7,x8,a1,a2,a3,a4,a5,a6,a7,a8,clk,ACC,p,out);
               input clk,p;
               input [24:0] x1,x2,x3,x4,x5,x6,x7,x8;
               input [63:0]a1,a2,a3,a4,a5,a6,a7,a8;
               output reg [63:0] ACC;
               output reg out;
               reg [31:0]i,c;
    reg [63:0]lout;
     reg [6:0]T;
     
     always@(posedge clk&p)
        begin 
        ACC=(-(a1+a2+a3+a4+a5+a6+a7+a8));
        ACC=({ACC[63],{63{1'b0}}})|(ACC>>1);
         i=0;c=0;  
       end
    
    always@(posedge clk&~p)
      begin  
       T[6]=(x1[i])^(x2[i]);
       T[5]=(x1[i])^(x3[i]);
       T[4]=(x1[i])^(x4[i]);
       T[3]=(x1[i])^(x5[i]);
       T[2]=(x1[i])^(x6[i]);
       T[1]=(x1[i])^(x7[i]);
       T[0]=(x1[i])^(x8[i]);
      i=i+1;
      lutout(a1,a2,a3,a4,a5,a6,a7,a8,T,lout);
      if(i<=24)  
          begin 
           if(~(x1[i-1]))
            begin
                ACC=ACC+lout;
                ACC=({ACC[63],{63{1'b0}}})|(ACC>>1);
                c=c+1;
              end
            else
            begin
                ACC=ACC-lout;
                ACC=({ACC[63],{63{1'b0}}})|(ACC>>1);
             end
           end
       else if(i==25)
       begin
           out=1;
           if((x1[i-1]))
                ACC=ACC+lout;
            else
                    ACC=ACC-lout;
           end
           else
           out=0;
      end
       task lutout;
           input [63:0]a1,a2,a3,a4,a5,a6,a7,a8;
           input [6:0]B;
           output reg [63:0]lout;
           reg [63:0] M1,
     M2  ,
     M3  ,
     M4  ,
     M5  ,
     M6  ,
     M7  ,
     M8  ,
     M9  ,
     M10 ,
     M11 ,
     M12 ,
     M13 ,
     M14 ,
     M15 ,
     M16 ,
     M17 ,
     M18 ,
     M19 ,
     M20 ,
     M21 ,
     M22 ,
     M23 ,
     M24 ,
     M25 ,
     M26 ,
     M27 ,
     M28 ,
     M29 ,
     M30 ,
     M31 ,
     M32 ,
     M33 ,
     M34 ,
     M35 ,
     M36 ,
     M37 ,
     M38 ,
     M39 ,
     M40 ,
     M41 ,
     M42 ,
     M43 ,
     M44 ,
     M45 ,
     M46 ,
     M47 ,
     M48 ,
     M49 ,
     M50 ,
     M51 ,
     M52 ,
     M53 ,
     M54 ,
     M55 ,
     M56 ,
     M57 ,
     M58 ,
     M59 ,
     M60 ,
     M61 ,
     M62 ,
     M63 ,
     M64 ,
     M65 ,
     M66 ,
     M67 ,
     M68 ,
     M69 ,
     M70 ,
     M71 ,
     M72 ,
     M73 ,
     M74 ,
     M75 ,
     M76 ,
     M77 ,
     M78 ,
     M79 ,
     M80 ,
     M81 ,
     M82 ,
     M83 ,
     M84 ,
     M85 ,
     M86 ,
     M87 ,
     M88 ,
     M89 ,
     M90 ,
     M91 ,
     M92 ,
     M93 ,
     M94 ,
     M95 ,
     M96 ,
     M97 ,
     M98 ,
     M99 ,
     M100,
     M101,
     M102,
     M103,
     M104,
     M105,
     M106,
     M107,
     M108,
     M109,
     M110,
     M111,
     M112,
     M113,
     M114,
     M115,
     M116,
     M117,
     M118,
     M119,
     M120,
     M121,
     M122,
     M123,
     M124,
     M125,
     M126,
     M127,M128;

           begin
M1  = (-(a1+a2+a3+a4+a5+a6+a7+a8));                           
M2  = (-(a1+a2+a3+a4+a5+a6+a7-a8));
M3  = (-(a1+a2+a3+a4+a5+a6-a7+a8));
M4  = (-(a1+a2+a3+a4+a5+a6-a7-a8));
M5  = (-(a1+a2+a3+a4+a5-a6+a7+a8));
M6  = (-(a1+a2+a3+a4+a5-a6+a7-a8));
M7  = (-(a1+a2+a3+a4+a5-a6-a7+a8));
M8  = (-(a1+a2+a3+a4+a5-a6-a7-a8));
M9  = (-(a1+a2+a3+a4-a5+a6+a7+a8));
M10  = (-(a1+a2+a3+a4-a5+a6+a7-a8));
M11  = (-(a1+a2+a3+a4-a5+a6-a7+a8));
M12  = (-(a1+a2+a3+a4-a5+a6-a7-a8));
M13  = (-(a1+a2+a3+a4-a5-a6+a7+a8));
M14  = (-(a1+a2+a3+a4-a5-a6+a7-a8));
M15  = (-(a1+a2+a3+a4-a5-a6-a7+a8));                                 
M16 = (-(a1+a2+a3+a4-a5-a6-a7-a8));
M17 = (-(a1+a2+a3-a4+a5+a6+a7+a8));
M18 = (-(a1+a2+a3-a4+a5+a6+a7-a8));
M19 = (-(a1+a2+a3-a4+a5+a6-a7+a8));
M20 = (-(a1+a2+a3-a4+a5+a6-a7-a8));
M21 = (-(a1+a2+a3-a4+a5-a6+a7+a8));
M22 = (-(a1+a2+a3-a4+a5-a6+a7-a8));
M23 =(- (a1+a2+a3-a4+a5-a6-a7+a8));
M24 = (-(a1+a2+a3-a4+a5-a6-a7-a8));
M25 = (-(a1+a2+a3-a4-a5+a6+a7+a8));
M26 = (-(a1+a2+a3-a4-a5+a6+a7-a8));
M27 = (-(a1+a2+a3-a4-a5+a6-a7+a8));
M28 = (-(a1+a2+a3-a4-a5+a6-a7-a8));
M29 = (-(a1+a2+a3-a4-a5-a6+a7+a8));
M30 = (-(a1+a2+a3-a4-a5-a6+a7-a8));
M31 = (-(a1+a2+a3-a4-a5-a6-a7+a8));
M32 = (-(a1+a2+a3-a4-a5-a6-a7-a8));
M33 = (-(a1+a2-a3+a4+a5+a6+a7+a8));
M34 = (-(a1+a2-a3+a4+a5+a6+a7-a8));
M35 = (-(a1+a2-a3+a4+a5+a6-a7+a8));
M36 = (-(a1+a2-a3+a4+a5+a6-a7-a8));
M37 = (-(a1+a2-a3+a4+a5-a6+a7+a8));
M38 = (-(a1+a2-a3+a4+a5-a6+a7-a8));
M39 = (-(a1+a2-a3+a4+a5-a6-a7+a8));
M40 = (-(a1+a2-a3+a4+a5-a6-a7-a8));
M41 = (-(a1+a2-a3+a4-a5+a6+a7+a8));
M42 = (-(a1+a2-a3+a4-a5+a6+a7-a8));
M43 = (-(a1+a2-a3+a4-a5+a6-a7+a8));
M44 = (-(a1+a2-a3+a4-a5+a6-a7-a8));
M45 = (-(a1+a2-a3+a4-a5-a6+a7+a8));
M46 = (-(a1+a2-a3+a4-a5-a6+a7-a8));
M47 = (-(a1+a2-a3+a4-a5-a6-a7+a8));
M48 = (-(a1+a2-a3+a4-a5-a6-a7-a8));
M49 = (-(a1+a2-a3-a4+a5+a6+a7+a8));
M50 = (-(a1+a2-a3-a4+a5+a6+a7-a8));
M51 = (-(a1+a2-a3-a4+a5+a6-a7+a8));
M52 = (-(a1+a2-a3-a4+a5+a6-a7-a8));
M53 = (-(a1+a2-a3-a4+a5-a6+a7+a8));
M54 = (-(a1+a2-a3-a4+a5-a6+a7-a8));
M55 = (-(a1+a2-a3-a4+a5-a6-a7+a8));
M56 = (-(a1+a2-a3-a4+a5-a6-a7-a8));
M57 = (-(a1+a2-a3-a4-a5+a6+a7+a8));
M58 = (-(a1+a2-a3-a4-a5+a6+a7-a8));
M59 = (-(a1+a2-a3-a4-a5+a6-a7+a8));
M60 = (-(a1+a2-a3-a4-a5+a6-a7-a8));
M61 = (-(a1+a2-a3-a4-a5-a6+a7+a8));
M62 = (-(a1+a2-a3-a4-a5-a6+a7-a8));
M63 = (-(a1+a2-a3-a4-a5-a6-a7+a8));
M64 = (-(a1+a2-a3-a4-a5-a6-a7-a8));
M65 = (-(a1-a2+a3+a4+a5+a6+a7+a8));
M66 = (-(a1-a2+a3+a4+a5+a6+a7-a8));
M67 = (-(a1-a2+a3+a4+a5+a6-a7+a8));
M68 = (-(a1-a2+a3+a4+a5+a6-a7-a8));
M69 = (-(a1-a2+a3+a4+a5+a6+a7+a8));
M70 = (-(a1-a2+a3+a4+a5-a6+a7-a8));
M71 = (-(a1-a2+a3+a4+a5-a6-a7+a8));
M72 = (-(a1-a2+a3+a4+a5-a6-a7-a8));
M73 = (-(a1-a2+a3+a4-a5+a6+a7+a8));
M74 = (-(a1-a2+a3+a4-a5+a6+a7-a8));
M75 = (-(a1-a2+a3+a4-a5+a6-a7+a8));
M76 = (-(a1-a2+a3+a4-a5+a6-a7-a8));
M77 = (-(a1-a2+a3+a4-a5-a6+a7+a8));
M78 = (-(a1-a2+a3+a4-a5-a6+a7-a8));
M79 = (-(a1-a2+a3+a4-a5-a6-a7+a8));
M80 = (-(a1-a2+a3+a4-a5-a6-a7-a8));
M81 = (-(a1-a2+a3-a4+a5+a6+a7+a8));
M82 = (-(a1-a2+a3-a4+a5+a6+a7-a8));
M83 = (-(a1-a2+a3-a4+a5+a6-a7+a8));
M84 = (-(a1-a2+a3-a4+a5+a6-a7-a8));
M85 = (-(a1-a2+a3-a4+a5-a6+a7+a8));
M86 = (-(a1-a2+a3-a4+a5-a6+a7-a8));
M87 = (-(a1-a2+a3-a4+a5-a6-a7+a8));
M88 = (-(a1-a2+a3-a4+a5-a6+a7-a8));
M89 = (-(a1-a2+a3-a4-a5+a6+a7+a8));
M90 = (-(a1-a2+a3-a4-a5+a6+a7-a8));
M91 = (-(a1-a2+a3-a4-a5+a6-a7+a8));
M92 = (-(a1-a2+a3-a4-a5+a6-a7-a8));
M93 = (-(a1-a2+a3-a4-a5-a6+a7+a8));
M94 = (-(a1-a2+a3-a4-a5-a6+a7-a8));
M95 = (-(a1-a2+a3-a4-a5-a6-a7+a8));
M96 = (-(a1-a2+a3-a4-a5-a6-a7-a8));
M97 = (-(a1-a2-a3+a4+a5+a6+a7+a8));
M98 = (-(a1-a2-a3+a4+a5+a6+a7-a8));
M99 = (-(a1-a2-a3+a4+a5+a6-a7+a8));
M100= (-(a1-a2-a3+a4+a5+a6-a7-a8));
M101= (-(a1-a2-a3+a4+a5-a6+a7+a8));
M102= (-(a1-a2-a3+a4+a5-a6+a7-a8));
M103= (-(a1-a2-a3+a4+a5-a6-a7+a8));
M104= (-(a1-a2-a3+a4+a5-a6-a7-a8));
M105= (-(a1-a2-a3+a4-a5+a6+a7+a8));
M106= (-(a1-a2-a3+a4-a5+a6+a7-a8));
M107= (-(a1-a2-a3+a4-a5+a6-a7+a8));
M108= (-(a1-a2-a3+a4-a5+a6-a7-a8));
M109= (-(a1-a2-a3+a4-a5-a6+a7+a8));
M110= (-(a1-a2-a3+a4-a5-a6+a7-a8));
M111= (-(a1-a2-a3+a4-a5-a6-a7+a8));
M112= (-(a1-a2-a3+a4-a5-a6-a7-a8));
M113= (-(a1-a2-a3-a4+a5+a6+a7+a8));
M114= (-(a1-a2-a3-a4+a5+a6+a7-a8));
M115= (-(a1-a2-a3-a4+a5+a6-a7+a8));
M116= (-(a1-a2-a3-a4+a5+a6-a7-a8));
M117= (-(a1-a2-a3-a4+a5-a6+a7+a8));
M118= (-(a1-a2-a3-a4+a5-a6+a7-a8));
M119= (-(a1-a2-a3-a4+a5-a6-a7+a8));
M120= (-(a1-a2-a3-a4+a5-a6-a7-a8));
M121= (-(a1-a2-a3-a4-a5+a6+a7+a8));
M122= (-(a1-a2-a3-a4-a5+a6+a7-a8));
M123= (-(a1-a2-a3-a4-a5+a6-a7+a8));
M124= (-(a1-a2-a3-a4-a5+a6-a7-a8));
M125= (-(a1-a2-a3-a4-a5-a6+a7+a8));
M126= (-(a1-a2-a3-a4-a5-a6+a7-a8));
M127= (-(a1-a2-a3-a4-a5-a6-a7+a8));
M128= (-(a1-a2-a3-a4-a5-a6-a7-a8));
     
case(B)
     0   :lout={M1[63],{63{1'b0}}} | (M1  >>1);
     1   :lout={M2[63],{63{1'b0}}} | (M2  >>1);
     2   :lout={M3[63],{63{1'b0}}} | (M3  >>1);
     3   :lout={M4[63],{63{1'b0}}} | (M4  >>1);
     4   :lout={M5[63],{63{1'b0}}} | (M5  >>1);
     5   :lout={M6[63],{63{1'b0}}} | (M6  >>1);
     6   :lout={M7[63],{63{1'b0}}} | (M7  >>1);
     7   :lout={M8[63],{63{1'b0}}} | (M8  >>1);
     8   :lout={M9[63],{63{1'b0}}} | (M9  >>1);
     9   :lout={M10[63],{63{1'b0}}} |(M10 >>1);
     10  :lout={M11[63],{63{1'b0}}} |(M11 >>1);
     11  :lout={M12[63],{63{1'b0}}} |(M12 >>1);
     12  :lout={M13[63],{63{1'b0}}} |(M13 >>1);
     13  :lout={M14[63],{63{1'b0}}} |(M14 >>1);
     14  :lout={M15[63],{63{1'b0}}} |(M15 >>1);
     15  :lout={M16[63],{63{1'b0}}} |(M16 >>1);
     16  :lout={M17[63],{63{1'b0}}} |(M17 >>1);
     17  :lout={M18[63],{63{1'b0}}} |(M18 >>1);
     18  :lout={M19[63],{63{1'b0}}} |(M19 >>1);
     19  :lout={M20[63],{63{1'b0}}} |(M20 >>1);
     20  :lout={M21[63],{63{1'b0}}} |(M21 >>1);
     21  :lout={M22[63],{63{1'b0}}} |(M22 >>1);
     22  :lout={M23[63],{63{1'b0}}} |(M23 >>1);
     23  :lout={M24[63],{63{1'b0}}} |(M24 >>1);
     24  :lout={M25[63],{63{1'b0}}} |(M25 >>1);
     25  :lout={M26[63],{63{1'b0}}} |(M26 >>1);
     26  :lout={M27[63],{63{1'b0}}} |(M27 >>1);
     27  :lout={M28[63],{63{1'b0}}} |(M28 >>1);
     28  :lout={M29[63],{63{1'b0}}} |(M29 >>1);
     29  :lout={M30[63],{63{1'b0}}} |(M30 >>1);
     30  :lout={M31[63],{63{1'b0}}} |(M31 >>1);
     31  :lout={M32[63],{63{1'b0}}} |(M32 >>1);
     32  :lout={M33[63],{63{1'b0}}} |(M33 >>1);
     33  :lout={M34[63],{63{1'b0}}} |(M34 >>1);
     34  :lout={M35[63],{63{1'b0}}} |(M35 >>1);
     35  :lout={M36[63],{63{1'b0}}} |(M36 >>1);
     36  :lout={M37[63],{63{1'b0}}} |(M37 >>1);
     37  :lout={M38[63],{63{1'b0}}} |(M38 >>1);
     38  :lout={M39[63],{63{1'b0}}} |(M39 >>1);
     39  :lout={M40[63],{63{1'b0}}} |(M40 >>1);
     40  :lout={M41[63],{63{1'b0}}} |(M41 >>1);
     41  :lout={M42[63],{63{1'b0}}} |(M42 >>1);
     42  :lout={M43[63],{63{1'b0}}} |(M43 >>1);
     43  :lout={M44[63],{63{1'b0}}} |(M44 >>1);
     44  :lout={M45[63],{63{1'b0}}} |(M45 >>1);
     45  :lout={M46[63],{63{1'b0}}} |(M46 >>1);
     46  :lout={M47[63],{63{1'b0}}} |(M47 >>1);
     47  :lout={M48[63],{63{1'b0}}} |(M48 >>1);
     48  :lout={M49[63],{63{1'b0}}} |(M49 >>1);
     49  :lout={M50[63],{63{1'b0}}} |(M50 >>1);
     50  :lout={M51[63],{63{1'b0}}} |(M51 >>1);
     51  :lout={M52[63],{63{1'b0}}} |(M52 >>1);
     52  :lout={M53[63],{63{1'b0}}} |(M53 >>1);
     53  :lout={M54[63],{63{1'b0}}} |(M54 >>1);
     54  :lout={M55[63],{63{1'b0}}} |(M55 >>1);
     55  :lout={M56[63],{63{1'b0}}} |(M56 >>1);
     56  :lout={M57[63],{63{1'b0}}} |(M57 >>1);
     57  :lout={M58[63],{63{1'b0}}} |(M58 >>1);
     58  :lout={M59[63],{63{1'b0}}} |(M59 >>1);
     59  :lout={M60[63],{63{1'b0}}} |(M60 >>1);
     60  :lout={M61[63],{63{1'b0}}} |(M61 >>1);
     61  :lout={M62[63],{63{1'b0}}} |(M62 >>1);
     62  :lout={M63[63],{63{1'b0}}} |(M63 >>1);
     63  :lout={M64[63],{63{1'b0}}} |(M64 >>1);
     64  :lout={M65[63],{63{1'b0}}} |(M65 >>1);
     65  :lout={M66[63],{63{1'b0}}} |(M66 >>1);
     66  :lout={M67[63],{63{1'b0}}} |(M67 >>1);
     67  :lout={M68[63],{63{1'b0}}} |(M68 >>1);
     68  :lout={M69[63],{63{1'b0}}} |(M69 >>1);
     69  :lout={M70[63],{63{1'b0}}} |(M70 >>1);
     70  :lout={M71[63],{63{1'b0}}} |(M71 >>1);
     71  :lout={M72[63],{63{1'b0}}} |(M72 >>1);
     72  :lout={M73[63],{63{1'b0}}} |(M73 >>1);
     73  :lout={M74[63],{63{1'b0}}} |(M74 >>1);
     74  :lout={M75[63],{63{1'b0}}} |(M75 >>1);
     75  :lout={M76[63],{63{1'b0}}} |(M76 >>1);
     76  :lout={M77[63],{63{1'b0}}} |(M77 >>1);
     77  :lout={M78[63],{63{1'b0}}} |(M78 >>1);
     78  :lout={M79[63],{63{1'b0}}} |(M79 >>1);
     79  :lout={M80[63],{63{1'b0}}} |(M80 >>1);
     80  :lout={M81[63],{63{1'b0}}} |(M81 >>1);
     81  :lout={M82[63],{63{1'b0}}} |(M82 >>1);
     82  :lout={M83[63],{63{1'b0}}} |(M83 >>1);
     83  :lout={M84[63],{63{1'b0}}} |(M84 >>1);
     84  :lout={M85[63],{63{1'b0}}} |(M85 >>1);
     85  :lout={M86[63],{63{1'b0}}} |(M86 >>1);
     86  :lout={M87[63],{63{1'b0}}} |(M87 >>1);
     87  :lout={M88[63],{63{1'b0}}} |(M88 >>1);
     88  :lout={M89[63],{63{1'b0}}} |(M89 >>1);
     89  :lout={M90[63],{63{1'b0}}} |(M90 >>1);
     90  :lout={M91[63],{63{1'b0}}} |(M91 >>1);
     91  :lout={M92[63],{63{1'b0}}} |(M92 >>1);
     92  :lout={M93[63],{63{1'b0}}} |(M93 >>1);
     93  :lout={M94[63],{63{1'b0}}} |(M94 >>1);
     94  :lout={M95[63],{63{1'b0}}} |(M95 >>1);
     95  :lout={M96[63],{63{1'b0}}} |(M96 >>1);
     96  :lout={M97[63],{63{1'b0}}} |(M97 >>1);
     97  :lout={M98[63],{63{1'b0}}} |(M98 >>1);
     98  :lout={M99[63],{63{1'b0}}} |(M99 >>1);
     99  :lout={M100[63],{63{1'b0}}} |(M100>>1);
     100 :lout={M101[63],{63{1'b0}}} |(M101>>1);
     101 :lout={M102[63],{63{1'b0}}} |(M102>>1);
     102 :lout={M103[63],{63{1'b0}}} |(M103>>1);
     103 :lout={M104[63],{63{1'b0}}} |(M104>>1);
     104 :lout={M105[63],{63{1'b0}}} |(M105>>1);
     105 :lout={M106[63],{63{1'b0}}} |(M106>>1);
     106 :lout={M107[63],{63{1'b0}}} |(M107>>1);
     107 :lout={M108[63],{63{1'b0}}} |(M108>>1);
     108 :lout={M109[63],{63{1'b0}}} |(M109>>1);
     109 :lout={M110[63],{63{1'b0}}} |(M110>>1);
     110 :lout={M111[63],{63{1'b0}}} |(M111>>1);
     111 :lout={M112[63],{63{1'b0}}} |(M112>>1);
     112 :lout={M113[63],{63{1'b0}}} |(M113>>1);
     113 :lout={M114[63],{63{1'b0}}} |(M114>>1);
     114 :lout={M115[63],{63{1'b0}}} |(M115>>1);
     115 :lout={M116[63],{63{1'b0}}} |(M116>>1);
     116 :lout={M117[63],{63{1'b0}}} |(M117>>1);
     117 :lout={M118[63],{63{1'b0}}} |(M118>>1);
     118 :lout={M119[63],{63{1'b0}}} |(M119>>1);
     119 :lout={M120[63],{63{1'b0}}} |(M120>>1);
     120 :lout={M121[63],{63{1'b0}}} |(M121>>1);
     121 :lout={M122[63],{63{1'b0}}} |(M122>>1);
     122 :lout={M123[63],{63{1'b0}}} |(M123>>1);
     123 :lout={M124[63],{63{1'b0}}} |(M124>>1);
     124 :lout={M125[63],{63{1'b0}}} |(M125>>1);
     125 :lout={M126[63],{63{1'b0}}} |(M126>>1);
     126 :lout={M127[63],{63{1'b0}}} |(M127>>1);
     127 :lout={M128[63],{63{1'b0}}} |(M128>>1);
     
             endcase
       end
       endtask              
endmodule